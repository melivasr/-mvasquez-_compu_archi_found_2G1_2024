module andOP(input logic [1:0] a,b, output logic [1:0] z);

assign z = a & b;

endmodule
